CircuitMaker Text
5.6
Probes: 2
Q1_2
Transient Analysis
0 247 502 65280
J2_2
Operating Point
0 279 386 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2030 58 2796 981
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
2198 154 2311 251
9961490 0
0
6 Title:
5 Name:
0
0
0
24
5 SIP3~
219 556 486 0 1 7
0 0
0
0 0 608 0
4 CONN
-13 -25 15 -17
5 IRRec
-14 -25 21 -17
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 J
4299 0 0
2
42116 0
0
5 SIP4~
219 552 623 0 1 9
0 0
0
0 0 608 0
4 CONN
9 2 37 10
5 RFRec
-17 -29 18 -21
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 J
9672 0 0
2
42116 0
0
5 SIP3~
219 212 285 0 1 7
0 0
0
0 0 608 180
4 CONN
-13 -25 15 -17
3 vr5
-13 -26 8 -18
0
0
0
0
0
3 vr5
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 J
7876 0 0
2
42116 0
0
5 SIP3~
219 193 193 0 1 7
0 0
0
0 0 608 180
4 CONN
-13 -25 15 -17
3 vr5
-13 -26 8 -18
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 J
6369 0 0
2
42116 0
0
5 SIP8~
219 134 450 0 8 17
0 19 20 21 14 22 23 24 25
0
0 0 608 180
4 CONN
9 2 37 10
2 J1
-13 -47 1 -39
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
1 J
9172 0 0
2
42116 0
0
5 SIP3~
219 53 279 0 3 7
0 9 26 2
0
0 0 608 0
4 CONN
-13 -25 15 -17
5 Screw
-14 -25 21 -17
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 J
7100 0 0
2
42116 1
0
5 SIP3~
219 104 279 0 3 7
0 9 5 2
0
0 0 608 0
4 CONN
-13 -25 15 -17
6 Switch
-19 -25 23 -17
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 J
3820 0 0
2
42116 2
0
5 SIP7~
219 65 377 0 7 15
0 27 28 29 30 31 2 5
0
0 0 608 0
4 CONN
-13 -43 15 -35
2 J4
-4 -43 10 -35
0
0
0
0
0
4 SIP7
15

0 1 2 3 4 5 6 7 1 2
3 4 5 6 7 0
0 0 0 512 1 0 0 0
1 J
7678 0 0
2
42116 3
0
5 SIP6~
219 68 453 0 6 13
0 32 33 34 35 36 37
0
0 0 608 0
4 CONN
9 2 37 10
2 J3
-7 -38 7 -30
0
0
0
0
0
4 SIP6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
0 0 0 512 1 0 0 0
1 J
961 0 0
2
42116 4
0
5 SIP6~
219 135 367 0 6 13
0 38 39 7 8 40 6
0
0 0 608 180
4 CONN
9 2 37 10
2 J2
-13 -38 1 -30
0
0
0
0
0
4 SIP6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
0 0 0 512 1 0 0 0
1 J
3178 0 0
2
42116 5
0
4 LED~
171 336 371 0 2 2
10 12 11
0
0 0 880 0
4 LED1
17 0 45 8
5 IRLED
14 -10 49 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3409 0 0
2
5.89705e-315 0
0
10 Capacitor~
219 446 517 0 2 5
0 13 2
0
0 0 832 90
5 .15uF
5 0 40 8
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3951 0 0
2
42116 6
0
4 LED~
171 107 591 0 2 2
10 10 2
0
0 0 880 0
4 LED1
17 0 45 8
4 YLED
17 -10 45 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8885 0 0
2
5.89705e-315 5.26354e-315
0
12 NPN Trans:C~
219 331 440 0 3 7
0 11 15 2
0
0 0 832 0
6 2N3904
18 0 60 8
2 Q2
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
81 0 0 0 1 0 0 0
1 Q
3780 0 0
2
5.89705e-315 5.30499e-315
0
7 Ground~
168 150 657 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
5.89705e-315 5.32571e-315
0
4 LED~
171 258 457 0 2 2
10 18 17
0
0 0 880 0
4 LED1
17 0 45 8
4 RLED
17 -10 45 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9442 0 0
2
42116 7
0
12 NPN Trans:C~
219 253 502 0 3 7
0 17 16 2
0
0 0 832 0
6 2N3904
18 0 60 8
2 Q1
32 -10 46 -2
0
0
14 %D %1 %2 %3 %M
0
0
4 SIP3
7

0 1 2 3 1 2 3 80425408
81 0 0 0 1 0 0 0
1 Q
9424 0 0
2
42116 8
0
9 Resistor~
219 107 556 0 2 5
0 10 8
0
0 0 864 90
3 330
7 0 28 8
2 R7
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
42116 9
0
9 Resistor~
219 352 572 0 4 5
0 6 2 0 -1
0
0 0 864 270
2 1M
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
42116 10
0
9 Resistor~
219 434 414 0 2 5
0 13 3
0
0 0 864 90
3 330
5 0 26 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
42116 11
0
9 Resistor~
219 336 336 0 2 5
0 12 4
0
0 0 864 90
2 56
7 0 21 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
5.89705e-315 5.38788e-315
0
9 Resistor~
219 209 440 0 2 5
0 14 15
0
0 0 864 0
3 330
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
5.89705e-315 5.39306e-315
0
9 Resistor~
219 211 502 0 2 5
0 14 16
0
0 0 864 0
3 330
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
5.89705e-315 5.39824e-315
0
9 Resistor~
219 258 414 0 2 5
0 18 4
0
0 0 864 90
2 56
7 0 21 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
42116 12
0
35
0 1 3 0 0 4224 0 0 2 21 0 5
409 203
409 604
515 604
515 610
540 610
2 0 4 0 0 4224 0 24 0 0 3 2
258 396
258 274
3 2 4 0 0 0 0 3 21 0 0 5
219 274
218 274
218 274
336 274
336 318
0 1 5 0 0 8192 0 0 3 17 0 4
166 312
166 320
219 320
219 292
2 0 2 0 0 12288 0 4 0 0 7 3
200 191
229 191
229 283
3 0 2 0 0 0 0 7 0 0 15 3
95 288
95 303
27 303
2 0 2 0 0 12288 0 3 0 0 15 4
219 283
229 283
229 325
27 325
0 0 2 0 0 0 0 0 0 32 24 2
148 611
258 611
2 0 2 0 0 0 0 12 0 0 27 2
446 508
446 487
2 0 2 0 0 0 0 19 0 0 27 2
352 590
352 611
1 6 6 0 0 8320 0 19 10 0 0 5
352 554
352 543
149 543
149 346
139 346
1 3 7 0 0 4224 0 1 10 0 0 6
547 477
225 477
225 463
166 463
166 373
139 373
2 4 8 0 0 8320 0 18 10 0 0 4
107 538
145 538
145 364
139 364
0 3 6 0 0 0 0 0 2 11 0 8
352 543
399 543
399 620
501 620
501 646
530 646
530 628
540 628
6 3 2 0 0 0 0 8 6 0 0 4
56 395
27 395
27 288
44 288
0 7 5 0 0 8320 0 0 8 17 0 4
86 312
44 312
44 404
56 404
2 1 5 0 0 0 0 7 4 0 0 8
95 279
83 279
83 312
166 312
166 241
208 241
208 200
200 200
1 1 9 0 0 12416 0 6 7 0 0 6
44 270
27 270
27 217
83 217
83 270
95 270
2 0 2 0 0 12416 0 13 0 0 15 4
107 601
107 609
28 609
28 395
1 1 10 0 0 4224 0 13 18 0 0 2
107 581
107 574
3 2 3 0 0 0 0 4 20 0 0 5
200 182
409 182
409 203
434 203
434 396
1 2 11 0 0 4224 0 14 11 0 0 2
336 422
336 381
1 1 12 0 0 4224 0 21 11 0 0 2
336 354
336 361
0 3 2 0 0 0 0 0 17 27 0 3
336 611
258 611
258 520
1 1 13 0 0 4224 0 20 12 0 0 4
434 432
434 537
446 537
446 526
1 3 13 0 0 16 0 12 1 0 0 5
446 526
446 537
502 537
502 495
547 495
2 3 2 0 0 0 0 1 14 0 0 7
547 486
446 486
446 487
428 487
428 611
336 611
336 458
4 0 2 0 0 0 0 2 0 0 27 6
540 637
540 654
487 654
487 627
384 627
384 611
1 0 14 0 0 8192 0 23 0 0 30 3
193 502
185 502
185 456
1 4 14 0 0 12416 0 22 5 0 0 4
191 440
185 440
185 456
138 456
2 2 15 0 0 4224 0 22 14 0 0 2
227 440
313 440
0 1 2 0 0 0 0 0 15 19 0 4
107 609
107 611
150 611
150 651
2 2 16 0 0 4224 0 23 17 0 0 2
229 502
235 502
2 1 17 0 0 4224 0 16 17 0 0 4
258 467
258 488
258 488
258 484
1 1 18 0 0 4224 0 24 16 0 0 2
258 432
258 447
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
