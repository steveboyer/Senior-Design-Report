CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
2030 58 2796 981
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
2198 154 2311 251
9961490 0
0
6 Title:
5 Name:
0
0
0
7
8 Antenna~
219 404 283 0 1 3
0 0
0
0 0 576 0
2 50
-8 -42 6 -34
4 ANT1
-14 -20 14 -12
0
0
10 %D %1 0 %V
0
0
3 BNC
3

0 1 1 0
82 0 0 0 0 0 0 0
3 ANT
5283 0 0
2
42116 0
0
5 SIP4~
219 378 362 0 1 9
0 0
0
0 0 608 0
4 CONN
9 2 37 10
7 RFtrans
-24 -29 25 -21
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
1 J
6874 0 0
2
42116 0
0
5 SIP3~
219 192 340 0 3 7
0 5 7 3
0
0 0 608 180
4 CONN
-13 -25 15 -17
5 Screw
-20 -26 15 -18
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 J
5305 0 0
2
5.89704e-315 0
0
5 SIP3~
219 193 385 0 3 7
0 2 8 4
0
0 0 608 180
4 CONN
-13 -25 15 -17
5 Screw
-20 -26 15 -18
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 1 0 0 0
1 J
34 0 0
2
5.89704e-315 0
0
7 Ground~
168 327 403 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
969 0 0
2
42116 0
0
4 LED~
171 327 293 0 2 2
10 6 2
0
0 0 880 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8402 0 0
2
5.89704e-315 0
0
9 Resistor~
219 327 250 0 2 5
0 6 3
0
0 0 864 90
3 330
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3751 0 0
2
5.89704e-315 5.30499e-315
0
8
1 1 0 0 0 0 0 2 1 0 0 5
366 349
340 349
340 317
404 317
404 299
0 1 2 0 0 8192 0 0 5 3 0 3
326 386
327 386
327 397
1 0 2 0 0 12416 0 4 0 0 8 5
200 392
211 392
211 386
327 386
327 376
3 2 3 0 0 16512 0 3 7 0 0 7
199 329
214 329
214 337
263 337
263 214
327 214
327 232
3 3 4 0 0 16528 0 4 2 0 0 5
200 374
200 377
242 377
242 367
366 367
1 2 5 0 0 16512 0 3 2 0 0 5
199 347
199 346
264 346
264 358
366 358
1 1 6 0 0 4224 0 7 6 0 0 2
327 268
327 283
2 4 2 0 0 0 0 6 2 0 0 3
327 303
327 376
366 376
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
